module conv5x5 (
    input clock,
    input reset,

    input [DWIDTH-1:0] data_in,
    input data_valid,

    output [DWIDTH-1:0] data_out,
    output data_valid_out

);
parameter DWIDTH = 8;

///
///

endmodule